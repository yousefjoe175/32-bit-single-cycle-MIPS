//MIPS module is the top module of the sytem which contains the interfacing
//between control unit, datapath unit, instruction memory, data memory
//it takes CLK and reset as input and test_value as an output 

module MIPS(
    input   wire            CLK,
    input   wire            reset,
    output  reg     [15:0]  test_value 
);



endmodule